# Language: Swedish (CP850)
# Translation courtesy of Martin Strömberg <ams@ludd.luth.se>.
# Needs translation for 1.13, 1.14, 1.15, 1.16, 1.17, 1.18, 2.12, 2.14, 2.15, 3.0, 3.1, 3.2, 3.3
#### Help        ####
1.0:Jämför två filer eller set av filer och visar skillnaderna mellan dem
1.1:FC [optioner] [drive1:][path1]filnamn1 [drive2][path2]filnamn2 [optioner]
1.2: /A    Visar bara den första och den sista raden för varje set av skillnader
1.3: /B    Gör en binär jämförelse
1.4: /C    Hantera gemener som versaler (problem med Å, Ä och Ö)
1.5: /L    Jämför filerna som ASCII-text.
1.6: /Mn   Sätt maximal antal skillnader vid binär jämförelse till n byte.
1.7:       (default = %d, 0 = ingen begränsning, /M = /M0)
1.8: /N    Visa radnumren vid textjämförelse
1.9: /S    Utöka jämförelsen till filerna i underkatalogerna
1.10: /T    Expandera inte tabbar till mellanslag
1.11: /W    Packa tabbar och mellanslag vid textjämförelse
1.12: /X    Visa inte kontextrader vid textjämförelse
1.13: /LBn  Set the maximum number of consecutive different ASCII lines to n
1.14: /nnn  Set the minimum number of consecutive matching lines to nnn
1.15:       for comparison resynchronization
1.16: /R    Show a brief final report (always active when using /S)
1.17: /Q    Don't show the list of differences
1.18: /U    Show the filenames of the files without a correspondent
#### Messages    ####
2.0:Ogiltig option: %s
2.1:För många filnamn
2.2:Ogiltigt filnamn
2.3:Ingen fil specifierad
2.4:Varning: filerna är olika stora!
2.5:Jämförelsen avslutad efter %d felträffar
2.6:Inga skillnader
2.7:Varning: jämförelsen avbruten efter %d rader
2.8:Otillräckligt med minne
2.9:Fel vid öppnande av fil %s
2.10:Jämför %s och %s
2.11:Ingen sådan fil eller katalog
2.12:Resync failed: files too different
2.13:Filerna är olika stora
2.14:The files are different
2.15:File %s has no correspondent (%s)
#### Report text ####
3.0:Compared %d files
3.1: in %d directories
3.2:%d files match, %d files are different
3.3:%d files have no correspondent
